`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.06.2025 19:40:53
// Design Name: 
// Module Name: Leading_Zero_Detector
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Leading_Zero_Detector(num,enable,count);
input [23:0]num;
input enable;
output reg [4:0]count;

always@(*) begin
    if(enable) begin
        casez (num)
        24'b1???????????????????????: count = 5'd0;
        24'b01??????????????????????: count = 5'd1;
        24'b001?????????????????????: count = 5'd2;
        24'b0001????????????????????: count = 5'd3;
        24'b00001???????????????????: count = 5'd4;
        24'b000001??????????????????: count = 5'd5;
        24'b0000001?????????????????: count = 5'd6;
        24'b00000001????????????????: count = 5'd7;
        24'b000000001???????????????: count = 5'd8;
        24'b0000000001??????????????: count = 5'd9;
        24'b00000000001?????????????: count = 5'd10;
        24'b000000000001????????????: count = 5'd11;
        24'b0000000000001???????????: count = 5'd12;
        24'b00000000000001??????????: count = 5'd13;
        24'b000000000000001?????????: count = 5'd14;
        24'b0000000000000001????????: count = 5'd15;
        24'b00000000000000001???????: count = 5'd16;
        24'b000000000000000001??????: count = 5'd17;
        24'b0000000000000000001?????: count = 5'd18;
        24'b00000000000000000001????: count = 5'd19;
        24'b000000000000000000001???: count = 5'd20;
        24'b0000000000000000000001??: count = 5'd21;
        24'b00000000000000000000001?: count = 5'd22;
        24'b000000000000000000000001: count = 5'd23;
        24'b000000000000000000000000: count = 5'd24;  // all zeros
        default: count = 5'd0;
    endcase
    end else begin
        count = 5'b0;
    end
end
endmodule
